# Translation by Martin Strömberg <ams@ludd.luth.se>.
0.0:Visa innehållet i en textfil en skärm i taget
0.1:Användning
0.2:kommando
0.3:fil
0.4:Tillgängliga tangenter
0.5:Nn
0.6:Nästa fil
0.7:Qq
0.8:Avsluta program
0.9:Mellanslag
0.10:Nästa sida
1.0:Okänd option
1.1:Ingen sådan fil
1.2:Kan inte öppna filen
2.0:Mera
2.1:<STDIN>
